	---------------------------------------------------------------------------------------------------
--
-- Title       : RNSsystem Compact RNS - extended Traditional
-- Design      : RNS systems
-- Author      : Gustavo Simas da Silva
-- Company     : SIPS INESC-id
--
---------------------------------------------------------------------------------------------------
--
-- File        : bin_adderTree.vhd
-- Generated   : Wed Oct  8 13:57:33 2012
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.20
--
---------------------------------------------------------------------------------------------------
--
-- Description : 
--
---------------------------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {CSA_2n_mp_1} architecture {Structural}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;   
--use work.bin_components.all;
--use work.compuRNS_def.all;
library work;
use work.fuctions.all;
--use work.rns_components.all;

entity LAB2b is
	generic (n : natural := 4);
	 port(SW   : in STD_LOGIC_VECTOR(4*n+1 downto 0);
			HEX1 : out STD_LOGIC_VECTOR(6 downto 0);
			HEX0 : out STD_LOGIC_VECTOR(6 downto 0));
end LAB2b;


--}} End of automatically maintained section

architecture Structural of LAB2b is

	component CSA_2n_mp_1 is
	generic (n : natural;
				-- modo = 0 => 2^n-1
				-- modo = 1 => 2^n+1
				modo: NATURAL);
  	 port(I0 : in STD_LOGIC_VECTOR((n-1) downto 0);
			I1 : in STD_LOGIC_VECTOR((n-1) downto 0);
			I2 : in STD_LOGIC_VECTOR((n-1) downto 0);
			S : out STD_LOGIC_VECTOR((n-1) downto 0);
			C : out STD_LOGIC_VECTOR((n-1) downto 0));
		end component;

  component adder_2n_mp_1 is 
	generic (n : natural :=4;
				-- modo = 0 => 2^n-1
				-- modo = 1 => 2^n+1
				modo: NATURAL := 0);
  	 port(A : in STD_LOGIC_VECTOR((n-1) downto 0);
			B : in STD_LOGIC_VECTOR((n-1) downto 0);
			S : out STD_LOGIC_VECTOR((n-1) downto 0);
			Cout: out STD_LOGIC);
	end component;
	
	component mux21 is
	generic (n : natural :=4);
	port (A: in std_logic_vector(n downto 0);
	B: in std_logic_vector(n downto 0);
	s: in std_logic;
	F: out std_logic_vector(n+1 downto 0)
	);
	end component;

  
  component Decod7seg is
	port (C: in std_logic_vector(3 downto 0);
	F: out std_logic_vector(6 downto 0)
	);
	end component;
  
signal zeros : std_logic_vector(n-1 downto 0);

signal cpa1_out: std_logic_vector(n downto 0);

signal cpa2_in1: std_logic_vector(n+1 downto 0);
signal cpa2_in2: std_logic_vector(n+1 downto 0);
signal cpa2_out: std_logic_vector(n+1 downto 0);

signal mux_out: std_logic_vector(n+1 downto 0);
signal disp1_sig: std_logic_vector(n-1 downto 0);

begin

converter : block

begin

cpa1: adder_2n_mp_1	generic map	(  n => n+1)
	                       port map ( A => SW(10 downto 6), B => SW(4 downto 0), S => cpa1_out);
							
csa1: CSA_2n_mp_1	generic map	(  n => n+2, modo => 0)
	                       port map ( I0 => SW(11 downto 6), I1 => SW(5 downto 0), I2 => SW(17 downto 12),
								  S => cpa2_in2, C => cpa2_in1);

cpa2: adder_2n_mp_1	generic map	(  n => n+2)
	                       port map ( A => cpa2_in1, B => cpa2_in2, S => cpa2_out);
								  
mux1: mux21	generic map	(  n => n)
	                       port map ( A => cpa2_out(4 downto 0), B => cpa1_out, s => cpa2_out(5), F => mux_out);

disp1_sig <= "00" & mux_out(5 downto 4);
								  
disp1: Decod7seg port map ( C => disp1_sig, F => HEX1);
disp2: Decod7seg port map ( C => mux_out(3 downto 0), F => HEX0);

end block;

end Structural;


